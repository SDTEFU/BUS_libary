// Generator : SpinalHDL v1.8.1    git head : 2a7592004363e5b40ec43e1f122ed8641cd8965b
// Component : SSM_BUS_test
// Git hash  : 4f05290e2b06b3d3417f1e984f0f1cb51ae029d4

`timescale 1ns/1ps

module SSM_BUS_test (
);



endmodule
